CONFIGURATION Fetch_PCVal_MUX_Fetch_PCVal_MUX_config OF Fetch_PCVal_MUX IS
   FOR Fetch_PCVal_MUX
   END FOR;
END Fetch_PCVal_MUX_Fetch_PCVal_MUX_config;