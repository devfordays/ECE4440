CONFIGURATION Mem_Multi16_Mem_Multi16_config OF Mem_Multi16 IS
   FOR Mem_Multi16
   END FOR;
END Mem_Multi16_Mem_Multi16_config;