--
-- VHDL Architecture Modic_Pipeline_lib.Multiplexor.Multiplexor
--
-- Created:
--          by - Owner.UNKNOWN (OWNER-PC)
--          at - 16:19:28 11/19/2012
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY Multiplexor IS
END ENTITY Multiplexor;

--
ARCHITECTURE Multiplexor OF Multiplexor IS
BEGIN
END ARCHITECTURE Multiplexor;

