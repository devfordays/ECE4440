CONFIGURATION Fetch_Mem_MUX_Fetch_Mem_MUX_config OF Fetch_Mem_MUX IS
   FOR Fetch_Mem_MUX
   END FOR;
END Fetch_Mem_MUX_Fetch_Mem_MUX_config;