CONFIGURATION Mem_Multi18_Mem_Multi18_config OF Mem_Multi18 IS
   FOR Mem_Multi18
   END FOR;
END Mem_Multi18_Mem_Multi18_config;