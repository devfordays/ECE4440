CONFIGURATION Decode_Right_MUX_Decode_Right_MUX_config OF Decode_Right_MUX IS
   FOR Decode_Right_MUX
   END FOR;
END Decode_Right_MUX_Decode_Right_MUX_config;