CONFIGURATION clock_clock_config OF clock IS
   FOR clock
   END FOR;
END clock_clock_config;