CONFIGURATION Reg_Reg_config OF Reg IS
   FOR Reg
   END FOR;
END Reg_Reg_config;