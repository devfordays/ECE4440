CONFIGURATION Fetch_PC_MUX_Fetch_PC_MUX_config OF Fetch_PC_MUX IS
   FOR Fetch_PC_MUX
   END FOR;
END Fetch_PC_MUX_Fetch_PC_MUX_config;