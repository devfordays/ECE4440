CONFIGURATION Execute_JumpUnit_Execute_JumpUnit_config OF Execute_JumpUnit IS
   FOR Execute_JumpUnit
   END FOR;
END Execute_JumpUnit_Execute_JumpUnit_config;