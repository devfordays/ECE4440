Modic_Pipeline_lib.Reg(Reg) :16:
Modic_Pipeline_lib.Reg(Reg) :4:
Modic_Pipeline_lib.Mem_Multi16(Mem_Multi16) rtlc_no_parameters
Modic_Pipeline_lib.Reg(Reg) :18:
Modic_Pipeline_lib.Mem_Multi1(Mem_Multi1) rtlc_no_parameters
Modic_Pipeline_lib.Register_Tracker_Control_MUX(Register_Tracker_Control_MUX) rtlc_no_parameters
Modic_Pipeline_lib.Register_File_four_sixteen_MUX(Register_File_four_sixteen_MUX) rtlc_no_parameters
Modic_Pipeline_lib.Register_File_TriState(Register_File_TriState) :16:
