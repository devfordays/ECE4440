--
-- VHDL Architecture Modic_Pipeline_lib.Top_Level_View.Top_Level_View
--
-- Created:
--          by - Owner.UNKNOWN (OWNER-PC)
--          at - 07:07:03 03/ 3/2013
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY Top_Level_View IS
-- Declarations

END Top_Level_View ;

--
ARCHITECTURE Top_Level_View OF Top_Level_View IS
BEGIN
END ARCHITECTURE Top_Level_View;

