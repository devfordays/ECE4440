-- Generation properties:
--   Format              : hierarchical
--   Generic mappings    : exclude
--   Leaf-level entities : direct binding
--   Regular libraries   : use library name
--   View name           : include
--   
CONFIGURATION tempor_struct_config OF tempor IS
   FOR struct
   END FOR;
END tempor_struct_config;
