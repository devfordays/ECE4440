CONFIGURATION Mem_new_MUX_Mem_new_MUX_config OF Mem_new_MUX IS
   FOR Mem_new_MUX
   END FOR;
END Mem_new_MUX_Mem_new_MUX_config;