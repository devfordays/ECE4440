CONFIGURATION Decode_MultSig_Decode_MultSig_config OF Decode_MultSig IS
   FOR Decode_MultSig
   END FOR;
END Decode_MultSig_Decode_MultSig_config;