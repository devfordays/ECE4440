CONFIGURATION Register_Tracker_Control_OR_Register_Tracker_Control_OR_config OF Register_Tracker_Control_OR IS
   FOR Register_Tracker_Control_OR
   END FOR;
END Register_Tracker_Control_OR_Register_Tracker_Control_OR_config;