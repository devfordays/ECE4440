CONFIGURATION Register_File_TriState_Register_File_TriState_config OF Register_File_TriState IS
   FOR Register_File_TriState
   END FOR;
END Register_File_TriState_Register_File_TriState_config;