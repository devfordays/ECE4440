CONFIGURATION Decode_Extra_MUX_Decode_Extra_MUX_config OF Decode_Extra_MUX IS
   FOR Decode_Extra_MUX
   END FOR;
END Decode_Extra_MUX_Decode_Extra_MUX_config;