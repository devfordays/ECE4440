CONFIGURATION Execute_Stage_ChangeNames_Execute_Stage_ChangeNames_config OF Execute_Stage_ChangeNames IS
   FOR Execute_Stage_ChangeNames
   END FOR;
END Execute_Stage_ChangeNames_Execute_Stage_ChangeNames_config;