--
-- VHDL Architecture Modic_Pipeline_lib.SRAM.SRAM
--
-- Created:
--          by - Owner.UNKNOWN (OWNER-PC)
--          at - 19:40:41 11/20/2012
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY SRAM IS
END ENTITY SRAM;

--
ARCHITECTURE SRAM OF SRAM IS
BEGIN
END ARCHITECTURE SRAM;

