CONFIGURATION Decode_Left_MUX_Decode_Left_MUX_config OF Decode_Left_MUX IS
   FOR Decode_Left_MUX
   END FOR;
END Decode_Left_MUX_Decode_Left_MUX_config;