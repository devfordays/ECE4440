CONFIGURATION Decode_Dest_MUX_Decode_Dest_MUX_config OF Decode_Dest_MUX IS
   FOR Decode_Dest_MUX
   END FOR;
END Decode_Dest_MUX_Decode_Dest_MUX_config;