CONFIGURATION Decode_Controller_Decode_Controller_config OF Decode_Controller IS
   FOR Decode_Controller
   END FOR;
END Decode_Controller_Decode_Controller_config;