CONFIGURATION Mem_Multiplexor_Mem_Multiplexor_config OF Mem_Multiplexor IS
   FOR Mem_Multiplexor
   END FOR;
END Mem_Multiplexor_Mem_Multiplexor_config;