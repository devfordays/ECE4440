CONFIGURATION Mem_Multi1_Mem_Multi1_config OF Mem_Multi1 IS
   FOR Mem_Multi1
   END FOR;
END Mem_Multi1_Mem_Multi1_config;