Modic_Pipeline_lib.Register_Tracker_Control_MUX(Register_Tracker_Control_MUX) rtlc_no_parameters
