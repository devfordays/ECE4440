CONFIGURATION easy_RAM_simu_behavior_config OF easy_RAM_simu IS
   FOR behavior
   END FOR;
END easy_RAM_simu_behavior_config;