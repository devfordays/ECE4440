Modic_Pipeline_lib.Mem_Multi16(Mem_Multi16) rtlc_no_parameters
Modic_Pipeline_lib.Mem_Multi1(Mem_Multi1) rtlc_no_parameters
