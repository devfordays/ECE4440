CONFIGURATION Fetch_Instr_MUX_Fetch_Instr_MUX_config OF Fetch_Instr_MUX IS
   FOR Fetch_Instr_MUX
   END FOR;
END Fetch_Instr_MUX_Fetch_Instr_MUX_config;