--
-- VHDL Architecture Modic_Pipeline_lib.james_code.james_code
--
-- Created:
--          by - Owner.UNKNOWN (OWNER-PC)
--          at - 15:33:43 03/ 3/2013
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY james_code IS
END ENTITY james_code;

--
ARCHITECTURE james_code OF james_code IS
BEGIN
END ARCHITECTURE james_code;

