--
-- VHDL Architecture Modic_Pipeline_lib.Instruction_StateMachine.Instruction_StateMachine
--
-- Created:
--          by - Owner.UNKNOWN (OWNER-PC)
--          at - 17:28:49 03/ 5/2013
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY Instruction_StateMachine IS
END ENTITY Instruction_StateMachine;

--
ARCHITECTURE Instruction_StateMachine OF Instruction_StateMachine IS
BEGIN
END ARCHITECTURE Instruction_StateMachine;

