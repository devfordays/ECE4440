CONFIGURATION Execute_ALU_Execute_ALU_config OF Execute_ALU IS
   FOR Execute_ALU
   END FOR;
END Execute_ALU_Execute_ALU_config;