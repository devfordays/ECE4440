CONFIGURATION Fetch_Incrementer_Fetch_Incrementer_config OF Fetch_Incrementer IS
   FOR Fetch_Incrementer
   END FOR;
END Fetch_Incrementer_Fetch_Incrementer_config;